package tta0_params is
  constant fu_LSU_dataw : integer := 32;
  constant fu_LSU_addrw : integer := 15;
end tta0_params;
